module spa
