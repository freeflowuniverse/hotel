module reception

struct Reception {

}

// Create Guest
// creates a new guest
fn (reception Reception) create_guest () {
	
}


