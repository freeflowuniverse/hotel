module vendor

pub interface IVendorClient {
	
}