module hr

// TODO is this redundant? is this what the employee supervisor is supposed to do?