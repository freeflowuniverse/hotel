module cleaning

// TODO clarify how this is structured