module actor_tests