module hoteldb