module flows

pub struct Vendor[T] {}

pub fn new_vendor[T]() {
	return Vendor[T]{}
}



