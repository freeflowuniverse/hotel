module accommodation

