module dock
