module department

// assuming that all requests are fairly similar
struct RequestHandlers {}

fn 