module flow_builder

/*
Given a Nodes struct:
- find the root flow
- 

*/