module restaurant