module hoteldb

pub struct Base{
pub mut:
	id string
	name string
	url string
	description string
	price string
	state ProductState	
}


//TODO: is there a way how to use our base?