module captain
