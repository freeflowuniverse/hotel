module cleaning

struct Cleaning {
	
}

// TODO clarify how this is structured