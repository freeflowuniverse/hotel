module flows

fn (flows ReceptionFlows)  (job ActionJob) {
	
}