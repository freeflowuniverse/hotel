module employee

import person

pub struct Employee {
	person.Person
}
