module telegram_bot

struct TelegramBot {
}