module spa

struct Spa {
	
}