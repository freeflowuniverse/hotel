module hotel


