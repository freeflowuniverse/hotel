module user


// import freeflowuniverse.baobab.jobs {ActionJob}
// import freeflowuniverse.hotel.actors.user

// fn (user IUser) get_user (identifier string, identifier_type string) !(IUser, string) {

// 	match identifier_type {
// 		'email' {
// 			if user.email == identifier { return user, user.type_name().all_after_last('.') }
// 		}
// 		'id' {
// 			if user.id == identifier { return user, user.type_name().all_after_last('.') }
// 		}
// 		'telegram_username' {
// 			if user.telegram_username == identifier { return user, user.type_name().all_after_last('.') }
// 		}
// 		else { return error("Invalid identifier type.")}
// 	}
// 	return error("Unrecognised identifier.")
// }	


