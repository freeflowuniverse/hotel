module main

import vweb
import os
import json

// ['/api/products'; get]
// ['/api/products/:id'; get]
// ['/api/products/strings'; get]
// ['/api/products/strings/:id'; get]