module vendor