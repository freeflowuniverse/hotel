module person

struct RequestHandlers {}

fn (rh RequestHandlers) function () ! {}