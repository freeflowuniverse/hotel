module cleaning
