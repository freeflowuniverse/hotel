module guest

import person

pub struct Guest {
	person.Person
}
