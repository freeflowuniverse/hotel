module actor_builder 

import os
import v.embed_file

pub struct SupervisorBuilder {
	actors []string
}

fn create_supervisor (actors []string, dir_path string) ! {
	
}