module vendor

pub struct VendorFlowsMixin {}